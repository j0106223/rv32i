module rv32_single_cycle_core (
    address,
    data,
);
    //instruction master
    //data master
endmodule